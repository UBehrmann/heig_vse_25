module regfile_assertions(
        input  logic      clk,
        input  logic[7:0] W,
        input  logic[7:0] A,
        input  logic[7:0] B,
        input  logic      Wen,
        input  logic[3:0] WA,
        input  logic[3:0] RAA,
        input  logic[3:0] RAB
);
endmodule
