-------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- Fichier      : packet_analyzer.vhd
--
-- Description  :
--
-- Auteur       : Yann Thoma
-- Date         : 07.10.2025
-- Version      : 0.1
--
-- Description  : Composant combinatoire pour l'analyse d'un paquet.
--
--| Modifications |------------------------------------------------------------
-- Version   Auteur Date               Description
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.packet_analyzer_pkg.all;

entity packet_analyzer is
    generic(
  		MAXSIZE : integer := 4;
        ERRNO : integer := 0
    );
    port(
        packet_i : in  std_logic_vector(MAXSIZE-1 downto 0);
        type_o   : out std_logic_vector(TYPESIZE-1 downto 0);
        length_o : out std_logic_vector(LENGTHSIZE-1 downto 0);
        error_o  : out std_logic_vector(ERRORSIZE-1 downto 0)
    );
end packet_analyzer;


`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
n5r4R7bodE3u7SMS6vDHRl+EcLIBmXhe4f+C9Mpy7X1Hkw4bys2oQ0pbwyzvCVIF
VA4IW/kapx9olSHX/Yi/Wpxi6h69M82wFtfECb921RjwozBYW4WNQsq5N3k0nplm
PKJSi7JZ8q84oJ4R2pKlJN1yz7KTuRHDMabkbho6toT+qQJV35YiRctK+ZSFwQW6
0c/iBSI5mlID0QcanFPrJPS3JKI3J6vIx7xtNNCbsZO60I7b2ivV9RvByHGZ1Z9M
+mQfyOehzQCTTS+XdLwCE/wDT5CZBkbf2s+bIAWM0pekN+2LaMDJunJJyMV4pfeY
jwlsXMc6PaZw6GfcRMHt0A==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7952 )
`protect data_block
WF3BaXwvFQJMqj0BCA03e0DwsEnxg2GlRAX3H/k9867uY8WrgN6UczQOWLacgRbT
ramcVNHYyQagr9JEA4ew09i2rfgutPYbQnGeNXrXESWCb2Lz2CP9NXqL6C0tNRz3
hhhUVSgt1hIpvfT/4m4rT8ZJa9uucXUfvx82QzXhs0gV3dN9idq9U4ekr2F7INkI
DiA1uXFBeHffSO+hY+yKwiucAe5Mi8ankw61JGv1Ib3lhqiNgQJ5SizHMZs1zjKS
Ur4fBtZSqOrOF253NuiNAnaS+joqQW52nlpmTQwFXsKtAzmJCeieerNQvxDLQ4G2
kwOFkPMkXoAEMzepxsgEJC22RO/ow1ebwMM5/V/ooU0oV3KlsdY5N1MAfc2iDdj7
cXrMphHxO2QkcbtSNe3fc9dKrFIZHxcv5Jrr9i57nUmSd+vY5Syd4uwMN4DuxB2r
bWVxt5uSdtNm0Tm173F97KRuSBXR9OYdwQ+CBiNlHBbz5q+bKlKjzziP/RMbEZPR
aZClNCRjnnGJNCP9A5bjkzQyaqCYa2jxFKDJ0a3C2ukCYtm3evi3LHK4ojA5rTUX
C3m1pjJZNpSA71CN79jXV4m2xCghqkad5xLVZNAmdy2TZyNu47/K61VGLza7YuYN
If1VyJwbxYEOGCAmIIUtkGNhpXIOn6nBLDYRt4uwehXA97WihbWnQWIzz+S6j3Jv
pbFWXe+jUAaihxucth4Sd87kry2uKbTDys3nZWn1tERzWCcL4r2vf0pZJFZgd6uh
P+5sHApguirAdrkUyEoc+bxRWy/vpRx1f71d+XXleJa20MAvriiBB+gxjmyyDnoh
rVO4dduv5qBVeAb2wivFldvGX//qyy7q6GvcarGov13ypFNSljnVlwdJiWFxxhpI
rnJ8vDxLaKeq/oC3eCYh+PTcTK9y6RTA4IjRWoBz2ggX+5WV6/xy7h3qyCTLz0Ra
zTrBPDcHVUlj00B2GpjsPjcoY1UMYbgMooociskMfoIPrWpTb0BXCgUnFQiO4kdW
jWYwZShG745oOBoxQKrNCKyTisrd0HEH/dhFKC/EiUQPxocP180BDHGaJcF3bCkM
l6AyZli/qNtYXy7ZWknYq56wvfkJVqpkFx1GFEhR7iMxqOOIAvAm3kLccl3qJ3e8
Zm6b0ehXsneV9Usyzp8iHj4rWKZfU9/GnnLQzhK5ttcVuIHkh7vuXPQDI3wosqMF
jH/6ALM2kduVfIuuLRm/6eRrDb7YZgcoDe1lUfBlt8Mo6Q3jdy77XzpZQ2awFXcl
tW5MOz78KEofxsQXsUafft8lN/Kzk9mh+DAHgzkjck6MRP5sr3bRNzAs07HfgZfW
Gju6l54G0xOGNS23jDX/Z+yxOXLVpzT6a3q5xnVUnY6lYctR0g+0n1lBWDPUTjfD
eCCDd16flbwBxlMaceJH6H4lrUpJIvWIMKKJAjISgzOfpZ2DFew95h3qf1Iq3Z1k
i73sfVmjE4ATL+U9WuLhMyXXuS1+AAuya4Vvx/BTsRSVBwHaoOD9UPValF08bw6r
mzkeYllLsUHE32mKLYnr45Ge8V4eb/7PmhOlSEVoD9gx9KKp+3YlC5xMZ72nWzRC
5ev7Y0J3aBEtRYx/AEEZTonnCh3tC1mVZH06NCVQh2F9ItUFWpUsRCkXtIV+/Z5d
RwkFnVzgHWZpN1c7gl9ACXjfcsVJ6ommAiW7F53y0YyoYBkJKsVTAUuZWugwfDf5
etk74ajQ9/umxTCDH/gxleMRwZuHmMC8thnFHvtzEQqoXlNYClb8RZs33iRgkVne
XDj+y/ANHBCyYi2FkZgZeMzvugbb0GPkiLjDS2k7nq5e8t4OG91Vh9IeN1vu53Nf
5Chj28jEc+Z2C11akj373IdbEcIcrjvHyMsG265XKBWx/u2edDRPmpQtrwYIiPWL
nf+In3J2ZGKV7jGGZuhMa4ipCxOwDaYA00Hplwsan02Qtl7iANNv25r5ptfDcmKA
LY/yollR2JtA+9Vf1IvHKngY3c1n5S7bOqXP5K6HCOlK1GZWMooKUOKpYjB4Lp1F
GBTU0d4atKXkzMBV/x4o3YqSIVJPTIp+Ujx7MLjzrNosl4S+47ZgQwAzhG6veNfo
ZYFRzbNjnYzKoJw7+0dTyKt5fjiq91F9C02JPqgCnl2g0brHb8+ZfyF+BFQ3z0DI
sG9GwgS+PE67CM0DFSvve73g3OD0WHxOk06DL5w1nGRr8qzISzUggn5PzrmMVXE/
0+eHgtWR+J5+jb2LRBg97/elVhyY9xXCjUlpor78QrfxYtShMKPIypJ5ROh8GYPD
xSX+d0b2wM3a7Rw/KFkfS5J3XJygHfeGaQwjMYVCS6FWURlYcnmOif/RuNgfpsNa
7UGucDeSe1oNyIHOd+jPjoO4hM8z1xGVphg1ZQOoJGXwYYUxf72CsJ4VfVzfXKoq
i4FJFuwqY515I4x9kN8nIojTx3zMVdwYoZB9rNxKxPj5ZKYNcx5qoHv5D/k3Gf/8
9mRxSaI/xO90d+Y6e+0z8btn/boqi0KsGAv2X24wFZx6e/Ukc4v0Vibp7XiwuNVo
/OlhYKZIirjKg7JQqmNTKHmYJjsZBkZPiK3+TRyGByColCFwK5DeLHwr2lVU3+4X
doX8QEerwDIFTgPZ93IkzpTPKwrtEaKi5wCGfQTnB87lFlBq2QjtAYivVT8XlcR7
SxStVhzwIFQCd8AofRC0KNJVloznQ13zPDSm5TZA0EW4a2o/f5e7K7o9Hdw7LZgv
zsz+2GMMTG52GgH1qDVC0Qm8YQwZGg3JhQG4v+nncxN+oKThxXz4NyJIzCF+4BLn
rb+pJQonoNS0Jkn7WRkSddoRWbA+8SefnPgSBQCI1CLShjPJzumxz862MCK0xaKS
tul3Qx+smnNz7usWGpWpxt0wsVfzFgBKYdhYoAccsrzwT2ZyhMUA+J0oLo/oNCOX
YtctoTyJI7FyHdht1z7+ADepPG5+wOmeAGGzm0jM8wFdz2jQ2/6B5nxu5VMWxjgy
1vsL6oynwex/gbAZRlLZcfu40qRu19MT17v58kwJZ7LnyU/0wd+Mg0YGlunKqtU/
YsTPpIccwz/7adKa4UIcsdmvDg4HoLLruy1b51ahUik1daqevi3zFjzFPE5f6wLT
400yyrSKq/2e7mTbiMsb+0CQn2hHVCFpe989C1ok9seUfDPJ9KgU9e4q9hVlV3/D
DO/nOrgIfYkmC6DPV2iTqGPahy5TvLgBzC8qJ4Fq6d+MsJZRkdYGzCAgNmRFw0KD
JXA8a5iBRcdgpsN+AcxETvJiB+jDuhfmGwS6zFemAiOV5F8bKPe+r/1wneJl37ho
AuL5nzNiFynmYCk8JxrcQ40S88dhgcrM+sKGleTCixt7VL4wQE8letwu8sSzL31e
FTNXCJSh6jeMTWmcftWg3Mzs3XrdKP4YD47uyr9CEPEF9/yOdUwTA9HYSDrd7PMt
meey7WkN1Sz+Ug4Dvsux1w7E8kH9jQZ81lLkTuDyv0HeuEtVQKose/Aq5ZedZTXw
n9TL5RRBnuGmDXowZVs2Vfnvy0gSX7eDRLvpSOoQpDkvlvJMwpDhDuY8OuJ2gi2p
l6Abq1xFx7iUGLF2YfUMdJZ8yCF0kp/Kj74ga4UAZGiPz76HWkZCmlMPgfPbMeNb
oRT9lYeKyQjwgAO/ZkxdDJnpTIEOH7tetdDRbotLEuC8QUXe55sthYz+5m60me7I
rN76wQaUiFDjWpq0L+9BAEmZnuyKlpAgTaoliCI+Otmv90NL6A68e0HQqyUXLXei
DjO9ZnUEc+OJOG/o/IZvXoYwhGroz262etVUesBP5Fsk9ZBmomoTF/eSrcqjZpl/
0VeAlol4rRcQiz754kuW88qZ38AijKKwyVod7DpvE+BbG4pTfJuA/GtMQTPg0VCt
pPrJDROlPSPgTNA5iPInK95rzMglXJKr/hQYg2OrOmoDoVvcGFDvtUlh5e1oJrTp
Y26xEsUi8BwCURY+JyewIjdQctfcl4RM4qQFQfHfugpTMvFYoECpU6JNynl6h6Ym
chiu8855erD2OvDdvcmeoILI8JbBalBfRtVzyKyL6lg6B4QgwddUTtOwUIYN0pw7
W4gqXU5m7hdqp26T4JuE4EZ3pg02Dw7piySwyK11Mp4eJMx1VUvUbvp8HFMG7C59
pdACZMY62ib5olW5auriBhQM2n3LtpqWWUj2cj4RNkkgX5+RUXvzxL9lZKjLaHOs
gCfHkfVEXRh97bx1PMSL1Vy8R2XW0yUPQRqFJPbALFawRMDMx+nAPbcWT1vU8a13
Cyj9Ecopp9bJFZianKaSmN0wGVz0OzbVGKki4vnurrxhTbIbYKCaAEyWD3COlScY
5WmfIDh9iAvsK6XcYYvl0tQcf6cB7BnMeOoNlGipnpYya3rz8AGuejXcPi5BQluM
rx+j9PAeznAC/Tx8ua7lSZsmDARErfw3cNrkpf4TdMYccXR664xvm0FN3jdrtDNe
qm0oZpoJNr/DHQeFZAdAkjwwliDdzUjFpF8rt+H1P6Jbdk+0Pl46GMCO81p8BSUL
5qydj9SBA8u7qzJO71Hpp4iHcUdnzTXPcZqKB5vhmImWyOGCH2pPkoIpvYiuSRLE
HQDd1t24WP5DIaoL87zq7E7zkVgZUna00VIUOGczk02BcG8dXNvSlXIx23Vu06Gz
lMMCGJvxWCIJ/2LdYYwRz8QxzJNWI2wXylgHDURicYHokvJgVaFs5jnE4OHKr8+5
1mLp13gtaOYZ/r6pIOJdqPWr4jHXHNAw/yLq07Xamc+9q84ydm56bLxZgBHJMcpU
bC9WBFKmX2DyI2pY0R9ykMfd13IX8c7AmjSoEUrgcroCLH1zqL+8sxUETxmf7fWn
4lQU0yuKGPgWPJXLK+rAsm3DBWMP/qB0BunA/8aJq3LFH2F93EhmVK4DiEbkF6NY
LH3tY5GQhc/r/hifhLahFpMgnqOl3CuOIoccVQCvW7L8sOrzkzeSXme1sxFYDvno
/7Ve5+EDqrjMMjAJVF6XXp8RzCO9xAV+iIW1EMFrZ36TWJiER6L19uFdbv0yw067
HhzqRMWcJG1mQffvJ8HdDoXBVl2lAWqx8vVhOHeqINiNAmUnuEzzXNmKabDv8qov
4xIZhxOKgapZIj9DBy0Y6c1kpm+Cbm2ulRkY/LOciR/uggzVhlCEfGx7JWc+BMPw
jWbNrnRhJ6vutE9XjnS5FGiu+5PDb+UtF9eOxk4rcGb/+FALAl0eRZSqqlA5XNwS
o2mqkeApM21RrfRLuLsoyVs+L2nZW2/WVgfooVZmlaUdQoiMpOYaboLUr6mTDhHC
PaqB+HknCnA9m+QwtbqEXfFFGKjH58RUL0ymJSKGnE30dIT7cWR6Qq4tnOMbrFr3
ctOdM5jFFhTgMnzL6M+GtPH4m+4c9ANCTneTiUIjYjiPEqw7f3mzVsU8I0Ow7TSh
zKI8+jLY3r/vUO3AB4ixX4o4EBoLdkEENMN/UVZP5z75CY00qOXrFy5b9Gw9dv0M
io+6XAUMVdV9MPYRmRxvqlToRMyK0SNAlF7pot3erOo6nxmGHXnmz1IrIyGrjEMm
t0lMPcDf4rymZFEU9BoNUb1DmkRfr4A5k+wkhVu2p3ZdM83vtYlJpUATbbu6VAKq
a83HFjGgBNjWAJsBMlUGwvEtNgBJI3Xh4lxO1gbxRwSDxNQvA18ZtFA3G3seLPN/
6em38vadnBRS3G3O7EeYJbd+8G3DKA9GkIgtA6T1kImHugXn1PjvAUlzonGiP3N1
OM1daKjX38PrpCBJqjwRzjQ3D0/9Gt+TOLtqY5LReaG9Ob7XEGw/UpGrRjgt6Bv1
QB+R64rwg0fmUkRplJLfE5P11S77FOgwLKwVoHNb0IAYwZ6HR9zb6kpNN7N10sne
lhBT5up15g0lKQINF696A+8IYouVAxHQULy9EmbhyONBh/IZ26jGbTVi/f1PvQ3R
8DCn/HjMu84AndIZKXaDo6/pYlx2B1HJdRGOfnPslw/R89QdEfxfnxj23VWJip1h
fZdzFsFwyDzlclrHNmLMNajZNgMtH5ohCXT80cPg1xZt9GcGZZ/MPq7AE5ErmaHL
vyaaEWgRN7nwtmWuYk3CT1L+pRYPYQ0PzDxON4o6CU8bUI+OAY9JienUpZZEDZQ/
EPV1qXkrRPHGGkvbnijHjAajBHUAnLcPIAdYqTzPnC586fP7pU9QmpWBVbQUpw0u
JmPKQ7NtQXTwdKYUCUXIcwAtd8hxlL4BEm88VaJ3sLNE6tUHxwzLc25tZnpOzTl3
bFKe4OlkUmAUcMY4cYgFVylFnSvLC/DGjNjGRacaini45cp5bVUrSVBfxKoAKSz0
9O9ML5fDaUFZvioUfGZWWjaLlKvSmPlLC9myc8G0QThXv7NxGWejfPIk2enUkJC6
Mk/iGzXqZFxYY2KTKfUjlY8MuvRLlO6vk4duYr+6ab0aLMt+cdulYYF0bNKONfRn
CPsW11XPPocie4uwEZGc+qxEMOzRlTYWTHwkR+3zUioHWoDNaaNTtlwMza5/feqR
kPjQ8WmuPcSv1Wt5h3YjfEHMP1HdxDwunPaA5mYnxWnfGLAM+dhYsuxj7E+83tNQ
CapZCzordKkw990UNXcPVyMJ16k+LbVLmCwRlXKhuUkrJvtMhuNdvyvM+e0LNI1e
NWPNjbh2Uon3Aimy89R6ya64vqATLcdoVw5Q5LHB42mjeZRa82hObkDOFCsUe4X+
Pwpk7lnUuiw85hBgBKJ39kiSzzWbrB3daWoV/8CpGz+uHH08eBOHVM7gk+EOk9/t
ti6Zf0Dhy5alUbR324tBBxTuRcBDwWtwhPZYGDN1yMS4Mu0j9K+GhSC3fa7Eyp2C
iMcxHmjTB25aHCICXfBwOi2xBpDR744fcSKfA6xmfebclId0tjvlWZWK1GsqYk79
UrJ1zUm0gAYf140l5g2YK8twcOAoJ9NY8e2xIbE2fs4voMNoNWmdPJrIyxS0k5oh
koi8bS3l7VBPVVl1w0EiVADOioWPfV/BLtrtfgIqXShTS5r/BKCVxXF2Owg2djWc
kSi7nSUH/9OTLSS9P42Kvuz26me2603/yYwdG2h1CursR0V8HTmiMGPUPn29ZK0G
aINl/FMpx6+F8GfxFhOYy8KoZMx0JVgqpzAoDhD1EaN8pCNIAUQPJOtKU70VVL72
x+qMnvEpIlH6r6xuO7mN6Wm1xo8/cBT8Di3wnNZXOOuOJ1OKVBYVHuQTq0RcKL0q
4AP735VmUgP32hVLKbKxkTTYOQ30ZoB4p4+3QadUtJthivciucuSjQJkFWplJ6Bf
lOumY8F676c7bNJNZxGrGyxDgnkVzLJ8C7SXIqt+3pNiP+7tnYY7XQztmZtKBoem
5TuRaKJdlyTERNQkD3V1QYkMqHMAJ7dH67+EuzgZIGWZWJZdClLQVB+00VokdfzA
xbVAoPgQ0STMXB4u+cyOTo4SP/udjLg7+ykzNA2M4jvtF3RbT25yWjn+drsj4LLE
E+TXbE+FgxE+MGhy8vWQDhlm/Sf0zlNm2inAGRNueX6BfZTKcIaWTWl/8aEZ5Lqa
MBHfYknB44FXZTx6AuPLCheIZs1ohziCfAP/W4Iqqe2aJBEJYc5YSZtLojRYLb79
XesjTQET7LSiPaANtMYiinKKm4v1LybuwAUiTGbQSv/yP6kD2bIxrgv9vvLzTSw8
BlcNlU8Lm8hLT41AgdpeWZRmKLe8NQAqBBb1uCWI/JD1hWh5emGOR5b4Mnx7rK+Y
dgjPTz7GRbAROlpVhJegCy2HNwrlFvlqx2pxyyqz56jWByzXBaxXhBLOIcVO+ivo
QicV7L5JntIMkOzmSneTeM85ERXLZCLdcvAvzQ8jDyphkL/AyvNcNb5UTQDv7x0P
GXOwHWgrOtjwi+PZOCuXToXLe0spr6+D2xb2Q948+4xFrftk8pERtsbVXVKS6oVT
hz3nar4G1SOTHbPTHGT3jJDvytiC7R9QHRqdew1lCEo6VY/hJlr3V6jBjK6OxNI9
t4e0OSNfHJ6de9i+NQygJDRIRDCt+Kpt4j92W8GcJyGitsmGMa1SoiUKZeHYKOpp
6nxoWx+/Hbev6hVBqP/jeiAQbHpTUj2xFuCH+QBsKyu+KH+M1p9rjZgsI5UgHry1
+FN8co948gI3yKXkuSHWt1fSLLEe37petAOJ20vcN+KMcjxTkkWAw+J4lKZPaSKb
itL77BqbVpDfxXBOFu7XMoc9LLuJhEcxBg1KNJa3qN+7M8wYrGacS9EBS11JEm/5
pHQtHih2qhA3q1ftRT33YEfDJMAO9cBW0oDK74u0VtFIXc2SYXgOAoHGfDvFoN/B
nYn4pEYqPXq4cwSBxjZ1nWk3Fx4lqoE7Yvku93TUTx5zR0L2Hszphu8T9SYluFIm
c5UwcQR7uUygzbmtoo4HAzxFqYjRIg2zuJbwVYHcprCcnpgj6K+fbQ7qENOspYz1
GhsLOepkBAozdefz/B2yEQac+YW4V3XqfNr2s477sxeaGJ5BSdudQ4y7E0W35vhM
qqkJf7FD5ixcIfNpuuoY5XfLSPE8beBorufh+9Q07TFfC1gnqRp+aw0ZwoXdLBSF
p1yaZc9J4EDYpy+nhEmwbhBAhOIX2WqTm9u6/ZIUUBwfAvY9L74jBTGA898UV6WY
6WIjTh3ltAxo/dOxvKU/lINKC+zquRic596u4dXefJO8NOuukZEC1r1pUyrK5X6T
GaBLlYnEAT2Fh0BAFbzuj7OScrs1Q+9lOVNxE1fZJA8e4e85OuzsewlhcN+Jn6jl
SwPlzoSuL61/Ckd5s7dX9KoxgHIB1ZHMOL7MMZYoL5H5SNr3WwX/7q47c0KIwK6I
Hi2nqnZspaFk3J/URyq7DKxB3yDpguaXQyUZ0aqh4KPxGHhabm8W270zb0ffmR5G
1+OvhESsJtnZDSFdcX+Y2DrkyA4AQPgzsOSW0CvqvM1yWhLIKUnLI+IF5vM9YaHI
Q3l6H8XKK7YlK1FvXZWtPGbT4QwMx0YhFOMxGkvVVI1H0WhD8DhDJCW/QWVUL1BH
zHVysW77/JFeQz0vMwfWzO7LpKYY3tkWAeya3jVkbWthsFP4iJwkfGUDx6gO9X/h
AQIUrnl/ePH0i/c6fjFMYpWsAOJ2wFU2WPhy4s3owE660uSHmCJCSwwTVVxz++/l
i7Kbb9YPPtB+c60/PKhCIVXIctf8JEoiEeJYwOMtkfoFZbVQRNjb8+dgsSHQ//1O
me9XHVwLOswjD240Gt7yrK6gNpeGRq/9jPmiaQfuYKZtQf4cvwSrhlfUyNxsT08K
rd006QB68kTKLeplipzMoLHosfSunFMow3KtC8HongYjwPXuhwMFzGfxxBCmovOt
0Fh13baErfhxW3oRfRqQPaI8UZsYH7Bj+woLpcNH9cV8KDxgAXTaPpMwApvbZKAM
Y1RPK+a76LBmwmQ5AfgwCIE83PXThL/MgDuIp5dwhoQ4LVfdFz22LWkIOGhprF1N
n7JwOhzqkmsLASt4wtT8T/Wr36KvI3nsBgy7OVm+mXkCFe9ex3WJQZ6YXfnog25X
h7KVZaWn0EsvzR4C2Gkze85/MhXIg+fO9ZwKQ8ap8xxjx3iw9f2I+Khnkvn09P7M
3CsjntCvWWd870At9/gkAHmk0gkkoN4bU8W6IjvXnxY9cXP8+eafqMrWvX5sVYgM
8ciNm+kZYyk42JBF3hBsRQaT3IveRTcInVeiYxI8LDl2hPZmEhrgSS62CYhz4C6/
qBwmE1D8Bbs8iGO/kodi0VB4De595mIvyuiBiM/PVLUjs5eaPOjp04bRF3mZJhF/
i436mqDpz4WYLzbXebL90odboP3zK5jOnnv4qKClQM1e+rdHuHctoRbH2l+zBIZ9
7WhIyvBF71C2iiTNiphoTNKTU5L3OWDhwCfxQHQvvtHCMqWSxu/u9v1pZYWcR3ZS
6vqqK5vG2+frTrBfXxNLyUKWItrgnAN6fmk45slECmUHx1HbAZBz6jOlYSjGJFs9
WXHJGuShdEh/7kR6ofs+TEE/ewVN+sDYokwU3UzFESins6QXbtacD7/W7Sb0X71I
QcReQt+VsERrna/xCnPslnRWXNgG02jpkVv/8r366mXRMPvi6OcUv8t/M8VFpdlW
sySlNwFtvOlQ76wj61uK3K9lOQfvtBM209jsucG7Tabw094pOuICC/MACKra4+H3
B+PhgkjIJCIFlcIgj/YC0KBvwR1kJn4ae5ldihSn/sB1m0LweqNA1izJxxXpzzSM
GTP/yrmnD2wv+G92VYfnjZI0xS5wNCanGLvVaTHQklbcgFINSkZE/wzHgmNIX3Lt
gT1qvVfnQZSRCmUnHwxbDundHR0lwcUYY8H64BVQxThk2T0MiSftLm3Ww4pMo4PD
B5v/UeCqilS7fS0KmzNBh9YRARGMgvnZVEyKyT2YUSry6SJhlzw/bJZ0rdOXwrC3
VEFOcs/xDxagj5SroSJLa4x2tFQSvIhGlIPK6RF5AJeR5xqF9oiJviM1gRzaPOTq
JUbXA7bQEnN9nHYoJuIebBoRJxQXBZ3YKlotaxmKX7TxcKRpty7nEPjLOuWoQzf8
UGXb8DO/a8QpTliiiMOYD5LncJkLiPmALBp/pUoKm0o=
`protect end_protected
